module pr_en (input [7:0] a,
              input [7:0] b,
              input [7:0] c,
              input [7:0] d,
              input [1:0] sel,
              output reg [7:0] out);

always @ (a or b or c or d or sel) begin
    if (sel == 2'b00)
        out <= a;
    else if (sel == 2'b01)
        out <= b;
    else if (sel == 2'b10)
        out <= c;
    else
        out <= d;
end
endmodule


module tb_4to1_mux;
    reg [7:0] a;
    reg [7:0] b;
    reg [7:0] c;
    reg [7:0] d;
    wire [7:0] out;
    reg [1:0] sel;
    integer i;
    
    pr_en    pr_en0 (.a (a),
    .b (b),
    .c (c),
    .d (d),
    .sel (sel),
    .out (out));
    
    initial begin
        $display(" == = TESTING PRIORITY ENCODER (4-to-1) CHIPVERIFY == = ");
        $monitor("Time = %0t: sel = %b, a = %b, b = %b, c = %b, d = %b", $time, sel, a, b, c, d);
        sel <= 0;
        a   <= $random;
        b   <= $random;
        c   <= $random;
        d   <= $random;
        
        for (i = 1; i < 4; i = i+1) begin
            #5 sel <= i;
        end
        
        #5 $finish;
    end
endmodule
