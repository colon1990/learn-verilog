module hello;
    initial
        begin
            $display("Hello world from haidh16: chip design class ");
            $finish;
        end
endmodule